module splitter (input [31:0] instruction,
	output reg [15:0] ,
	output reg [] address;
	output reg [4:0] rs,
	output reg [4:0] rt,
	output reg [4:0] rd,
	output reg [5:0] op,
	output reg [5:0] func);

always @(*) begin

end
endmodule
