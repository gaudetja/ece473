module splitter (input [31:0] instruction,
	output reg [15:0] offset,
	output reg [4:0] rs,
	output reg [4:0] rt,
	output reg [4:0] rd,
	output reg [5:0] op);

always @(*) begin

end
endmodule
