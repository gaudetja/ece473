module controller(input [6:0] op, output reg [2:0] alucontrol, output reg [5:0] muxout);
always @(*)
begin

end
endmodule
