//Add two 8bit numbers without carry


module plusfour (input [31:0] INPUT, output [31:0] SUM);

assign SUM = INPUT + 4;

endmodule
