//Add two 8bit numbers without carry


module plusfour (input [7:0] INPUT, output [7:0] SUM);

assign SUM = INPUT + 4;

endmodule
