//Add two 8bit numbers without carry


module bitadder (input [7:0] NUMBER1, input [7:0] NUMBER2, output [7:0] SUM);

assign SUM = NUMBER1 + NUMBER2;

endmodule
